`include "src/CSA.v"

module tb;

    module CSA_Adder32 ();

    
    
endmodule